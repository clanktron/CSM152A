module stopwatch(SEL, ADJ);

    input [7:0] SEL, ADJ;

    always
