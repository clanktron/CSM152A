module counter(SEL, ADJ, RESET, PAUSE, onehz, twohz, speedyhz, blinkyhz);

    input SEL, ADJ;

    always

