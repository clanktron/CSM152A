module stopwatch(SEL, ADJ, RESET, PAUSE);

    input SEL, ADJ, RESET, PAUSE;

    always @ (posedge clk) begin

    end
